module interrupt_controller